`timescale 1ns/1ps

module testbench();

    reg [3:0]IN;
    wire odd_out,even_out;

    four_bit_PARITY_always fbfal (
      .IN(IN),
      .odd_out(odd_out),
      .even_out(even_out)
    );

    initial
    begin
        IN = 4'b0000;
        #10 IN = 4'b0001;
        #10 IN = 4'b0010;
        #10 IN = 4'b0011;
        #10 IN = 4'b0100;
        #10 IN = 4'b0101;
        #10 IN = 4'b0110;
        #10 IN = 4'b0111;
        
        #10 IN = 4'b1000;
        #10 IN = 4'b1001;
        #10 IN = 4'b1010;
        #10 IN = 4'b1011;
        #10 IN = 4'b1100;
        #10 IN = 4'b1101;
        #10 IN = 4'b1110;
        #10 IN = 4'b1111;
        #10 ;

    end

endmodule