// 모듈

// 모듈 : Verilog에서 기본적인 설계 블록이다. 모듈은 요소 또는 하위 수준 설계 블록의 집합이다.
// 일반적으로 요소는 설계시 자주 사용되는 공통의 기능을 제공하기 위해 그룹지어서 모듈에 포함된다.
// 모듈은 포트 인터페이스를 통해서 상위 수준의 블록에 필요한 기능을 제공해주지만, 내부 구현은 숨긴다.
// 이것은 설계자가 다은 부분에 영향을 주지 않고 모듈의 내부를 수정할 수 있게 해준다.


// 모듈 예
module <모듈 이름>(<모듈 터미널 리스트>);
...
< 모듈 내용 >
...
...
endmodule


//=> T_FF 모듈 정의
module T_FF(q,clock,reset);
.
.
< T-FF기능>
.
.
endmodule


// Verilog는 행위적이고 구조적인 언어이다.
// 각 모듈의 내부는 설계의 쓰임에 따라 4가지 추상화 수준으로 정의할 수있다.
// 모듈은 추상화 수준과 관계없이 외부에서는 갗게 동작한다.
// 모듈의 내부는 외부로부터 숨겨져 있다.

// 행위 또는 알고리즘 수준(Behavioral or algorithmic level)
// Verilog에서 제공하는 추상화의 가장 상위 수준이다.
// 자세한 하드웨어구현에 관계없이 원하는 디자인 알고리즘을 바로 사용함으로써 모듈을 구현한다.

// 데이터플로우 수준(Dataflow level)
// 데이터의 흐름을 명백히 나타냄으로써 모듈을 구현한다. 
// 설계자는 하드웨어 레지스터 사이의 데이터 흐름과 데이터가 어떨게 처리되는지를 알고 있어야한다.

// 게이트 수준(Switch level)
// 논리 게이트와 게이트 사이의 연결에 의해 모듈이 구현된다.
// 이 수준에서의 설계는 게이트 수준 논리 다이어그램에 의해 묘사하는 것과 유사하다.

// 스위치 수준(Switch level)
// Verilog에서 제공하는 추상화의 가장 하위 수준이다.
// 스위치와 기억노드, 그리고 그것들의 연결에 의해서 모듈이 구현된다.


// 디지털 설계에서 레지스터 전송 수준(RTL)이라는 용어는
// 종종 행위 수준구조와 데이터 플로우수준 구조를 썩어서 사용하는 Verilog표현을 뜻하고
// 이는 논리 합성 도구의 입력으로 사용 가능하다.